`include "uvm_macros.svh"
import uvm_pkg::*;
//`include "apb_design.sv"

`include "defines.svh"
`include "ApbInterface.sv"
`include "ApbSeqItem.sv"
`include "ApbSequence.sv"
`include "ApbSequencer.sv"
`include "ApbDriver.sv"
`include "ApbIpMonitor.sv"
`include "ApbOpMonitor.sv"
`include "ApbActiveAgent.sv"
`include "ApbPassiveAgent.sv"
`include "ApbScoreboard.sv"
`include "ApbCoverage.sv"
`include "ApbEnvironment.sv"
`include "ApbTest.sv"

