`define AW 9
`define DW 9
